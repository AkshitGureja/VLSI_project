magic
tech scmos
timestamp 1638853031
<< nwell >>
rect -20 3 311 23
rect -20 -50 319 -30
rect 225 -51 319 -50
rect -20 -103 297 -83
rect -20 -156 308 -136
<< ntransistor >>
rect -9 -15 -7 -11
rect 3 -15 5 -11
rect 19 -15 21 -11
rect 38 -15 40 -11
rect 54 -15 56 -11
rect 70 -15 72 -11
rect 86 -15 88 -11
rect 102 -15 104 -11
rect 118 -15 120 -11
rect 134 -15 136 -11
rect 144 -15 146 -11
rect 160 -15 162 -11
rect 176 -15 178 -11
rect 186 -15 188 -11
rect 202 -15 204 -11
rect 218 -15 220 -11
rect 234 -15 236 -11
rect 250 -15 252 -11
rect 266 -15 268 -11
rect 282 -15 284 -11
rect 298 -15 300 -11
rect -9 -68 -7 -64
rect 3 -68 5 -64
rect 19 -68 21 -64
rect 38 -68 40 -64
rect 54 -68 56 -64
rect 70 -68 72 -64
rect 86 -68 88 -64
rect 94 -68 96 -64
rect 104 -68 106 -64
rect 120 -68 122 -64
rect 136 -68 138 -64
rect 146 -68 148 -64
rect 162 -68 164 -64
rect 178 -68 180 -64
rect 186 -68 188 -64
rect 194 -68 196 -64
rect 210 -68 212 -64
rect 226 -68 228 -64
rect 234 -68 236 -64
rect 242 -68 244 -64
rect 258 -68 260 -64
rect 274 -68 276 -64
rect 290 -68 292 -64
rect 306 -68 308 -64
rect -9 -121 -7 -117
rect 3 -121 5 -117
rect 19 -121 21 -117
rect 38 -121 40 -117
rect 54 -121 56 -117
rect 70 -121 72 -117
rect 86 -121 88 -117
rect 94 -121 96 -117
rect 102 -121 104 -117
rect 112 -121 114 -117
rect 128 -121 130 -117
rect 144 -121 146 -117
rect 152 -121 154 -117
rect 160 -121 162 -117
rect 168 -121 170 -117
rect 184 -121 186 -117
rect 200 -121 202 -117
rect 209 -121 211 -117
rect 225 -121 227 -117
rect 241 -121 243 -117
rect 251 -121 253 -117
rect 259 -121 261 -117
rect 267 -121 269 -117
rect 283 -121 285 -117
rect -9 -174 -7 -170
rect 3 -174 5 -170
rect 19 -174 21 -170
rect 38 -174 40 -170
rect 54 -174 56 -170
rect 70 -174 72 -170
rect 86 -174 88 -170
rect 94 -174 96 -170
rect 102 -174 104 -170
rect 110 -174 112 -170
rect 120 -174 122 -170
rect 136 -174 138 -170
rect 152 -174 154 -170
rect 161 -174 163 -170
rect 169 -174 171 -170
rect 185 -174 187 -170
rect 201 -174 203 -170
rect 210 -174 212 -170
rect 226 -174 228 -170
rect 242 -174 244 -170
rect 250 -174 252 -170
rect 259 -174 261 -170
rect 268 -174 270 -170
rect 277 -174 279 -170
rect 295 -174 297 -170
<< ptransistor >>
rect -9 9 -7 17
rect 3 9 5 17
rect 19 9 21 17
rect 38 9 40 17
rect 54 9 56 17
rect 70 9 72 17
rect 86 9 88 17
rect 102 9 104 17
rect 118 9 120 17
rect 134 9 136 17
rect 144 9 146 17
rect 160 9 162 17
rect 176 9 178 17
rect 186 9 188 17
rect 202 9 204 17
rect 218 9 220 17
rect 234 9 236 17
rect 250 9 252 17
rect 266 9 268 17
rect 282 9 284 17
rect 298 9 300 17
rect -9 -44 -7 -36
rect 3 -44 5 -36
rect 19 -44 21 -36
rect 38 -44 40 -36
rect 54 -44 56 -36
rect 70 -44 72 -36
rect 86 -44 88 -36
rect 94 -44 96 -36
rect 104 -44 106 -36
rect 120 -44 122 -36
rect 136 -44 138 -36
rect 146 -44 148 -36
rect 162 -44 164 -36
rect 178 -44 180 -36
rect 186 -44 188 -36
rect 194 -44 196 -36
rect 210 -44 212 -36
rect 226 -44 228 -36
rect 234 -44 236 -36
rect 242 -44 244 -36
rect 258 -44 260 -36
rect 274 -44 276 -36
rect 290 -44 292 -36
rect 306 -44 308 -36
rect -9 -97 -7 -89
rect 3 -97 5 -89
rect 19 -97 21 -89
rect 38 -97 40 -89
rect 54 -97 56 -89
rect 70 -97 72 -89
rect 86 -97 88 -89
rect 94 -97 96 -89
rect 102 -97 104 -89
rect 112 -97 114 -89
rect 128 -97 130 -89
rect 144 -97 146 -89
rect 152 -97 154 -89
rect 160 -97 162 -89
rect 168 -97 170 -89
rect 184 -97 186 -89
rect 200 -97 202 -89
rect 209 -97 211 -89
rect 225 -97 227 -89
rect 241 -97 243 -89
rect 251 -97 253 -89
rect 259 -97 261 -89
rect 267 -97 269 -89
rect 283 -97 285 -89
rect -9 -150 -7 -142
rect 3 -150 5 -142
rect 19 -150 21 -142
rect 38 -150 40 -142
rect 54 -150 56 -142
rect 70 -150 72 -142
rect 86 -150 88 -142
rect 94 -150 96 -142
rect 102 -150 104 -142
rect 110 -150 112 -142
rect 120 -150 122 -142
rect 136 -150 138 -142
rect 152 -150 154 -142
rect 161 -150 163 -142
rect 169 -150 171 -142
rect 185 -150 187 -142
rect 201 -150 203 -142
rect 210 -150 212 -142
rect 226 -150 228 -142
rect 242 -150 244 -142
rect 250 -150 252 -142
rect 259 -150 261 -142
rect 268 -150 270 -142
rect 277 -150 279 -142
rect 295 -150 297 -142
<< ndiffusion >>
rect -10 -15 -9 -11
rect -7 -15 3 -11
rect 5 -15 6 -11
rect 18 -15 19 -11
rect 21 -15 22 -11
rect 37 -15 38 -11
rect 40 -15 41 -11
rect 45 -15 49 -11
rect 53 -15 54 -11
rect 56 -15 57 -11
rect 69 -15 70 -11
rect 72 -15 73 -11
rect 85 -15 86 -11
rect 88 -15 89 -11
rect 93 -15 97 -11
rect 101 -15 102 -11
rect 104 -15 105 -11
rect 117 -15 118 -11
rect 120 -15 121 -11
rect 133 -15 134 -11
rect 136 -15 144 -11
rect 146 -15 147 -11
rect 159 -15 160 -11
rect 162 -15 163 -11
rect 175 -15 176 -11
rect 178 -15 180 -11
rect 184 -15 186 -11
rect 188 -15 189 -11
rect 201 -15 202 -11
rect 204 -15 205 -11
rect 217 -15 218 -11
rect 220 -15 221 -11
rect 225 -15 229 -11
rect 233 -15 234 -11
rect 236 -15 237 -11
rect 249 -15 250 -11
rect 252 -15 253 -11
rect 265 -15 266 -11
rect 268 -15 269 -11
rect 273 -15 277 -11
rect 281 -15 282 -11
rect 284 -15 285 -11
rect 297 -15 298 -11
rect 300 -15 301 -11
rect -10 -68 -9 -64
rect -7 -68 3 -64
rect 5 -68 6 -64
rect 18 -68 19 -64
rect 21 -68 22 -64
rect 37 -68 38 -64
rect 40 -68 41 -64
rect 45 -68 49 -64
rect 53 -68 54 -64
rect 56 -68 57 -64
rect 69 -68 70 -64
rect 72 -68 73 -64
rect 85 -68 86 -64
rect 88 -68 94 -64
rect 96 -68 104 -64
rect 106 -68 107 -64
rect 119 -68 120 -64
rect 122 -68 123 -64
rect 135 -68 136 -64
rect 138 -68 146 -64
rect 148 -68 149 -64
rect 161 -68 162 -64
rect 164 -68 165 -64
rect 177 -68 178 -64
rect 180 -68 186 -64
rect 188 -68 194 -64
rect 196 -68 197 -64
rect 209 -68 210 -64
rect 212 -68 213 -64
rect 225 -68 226 -64
rect 228 -68 229 -64
rect 233 -68 234 -64
rect 236 -68 237 -64
rect 241 -68 242 -64
rect 244 -68 245 -64
rect 257 -68 258 -64
rect 260 -68 261 -64
rect 273 -68 274 -64
rect 276 -68 277 -64
rect 281 -68 285 -64
rect 289 -68 290 -64
rect 292 -68 293 -64
rect 305 -68 306 -64
rect 308 -68 309 -64
rect -10 -121 -9 -117
rect -7 -121 3 -117
rect 5 -121 6 -117
rect 18 -121 19 -117
rect 21 -121 22 -117
rect 37 -121 38 -117
rect 40 -121 41 -117
rect 45 -121 49 -117
rect 53 -121 54 -117
rect 56 -121 57 -117
rect 69 -121 70 -117
rect 72 -121 73 -117
rect 85 -121 86 -117
rect 88 -121 94 -117
rect 96 -121 102 -117
rect 104 -121 112 -117
rect 114 -121 115 -117
rect 127 -121 128 -117
rect 130 -121 131 -117
rect 143 -121 144 -117
rect 146 -121 152 -117
rect 154 -121 160 -117
rect 162 -121 168 -117
rect 170 -121 171 -117
rect 183 -121 184 -117
rect 186 -121 187 -117
rect 199 -121 200 -117
rect 202 -121 209 -117
rect 211 -121 212 -117
rect 224 -121 225 -117
rect 227 -121 228 -117
rect 240 -121 241 -117
rect 243 -121 244 -117
rect 248 -121 251 -117
rect 253 -121 254 -117
rect 258 -121 259 -117
rect 261 -121 262 -117
rect 266 -121 267 -117
rect 269 -121 270 -117
rect 282 -121 283 -117
rect 285 -121 286 -117
rect -10 -174 -9 -170
rect -7 -174 3 -170
rect 5 -174 6 -170
rect 18 -174 19 -170
rect 21 -174 22 -170
rect 37 -174 38 -170
rect 40 -174 41 -170
rect 45 -174 49 -170
rect 53 -174 54 -170
rect 56 -174 57 -170
rect 69 -174 70 -170
rect 72 -174 73 -170
rect 85 -174 86 -170
rect 88 -174 94 -170
rect 96 -174 102 -170
rect 104 -174 110 -170
rect 112 -174 120 -170
rect 122 -174 123 -170
rect 135 -174 136 -170
rect 138 -174 139 -170
rect 151 -174 152 -170
rect 154 -174 161 -170
rect 163 -174 169 -170
rect 171 -174 172 -170
rect 184 -174 185 -170
rect 187 -174 188 -170
rect 200 -174 201 -170
rect 203 -174 210 -170
rect 212 -174 213 -170
rect 225 -174 226 -170
rect 228 -174 229 -170
rect 241 -174 242 -170
rect 244 -174 245 -170
rect 249 -174 250 -170
rect 252 -174 254 -170
rect 258 -174 259 -170
rect 261 -174 263 -170
rect 267 -174 268 -170
rect 270 -174 271 -170
rect 275 -174 277 -170
rect 279 -174 282 -170
rect 294 -174 295 -170
rect 297 -174 298 -170
<< pdiffusion >>
rect -10 9 -9 17
rect -7 9 -4 17
rect 0 9 3 17
rect 5 9 6 17
rect 18 9 19 17
rect 21 9 22 17
rect 37 9 38 17
rect 40 9 41 17
rect 53 9 54 17
rect 56 9 57 17
rect 69 9 70 17
rect 72 9 73 17
rect 85 9 86 17
rect 88 9 89 17
rect 101 9 102 17
rect 104 9 105 17
rect 117 9 118 17
rect 120 9 121 17
rect 133 9 134 17
rect 136 9 138 17
rect 142 9 144 17
rect 146 9 147 17
rect 159 9 160 17
rect 162 9 163 17
rect 175 9 176 17
rect 178 9 186 17
rect 188 9 189 17
rect 201 9 202 17
rect 204 9 205 17
rect 217 9 218 17
rect 220 9 221 17
rect 233 9 234 17
rect 236 9 237 17
rect 249 9 250 17
rect 252 9 253 17
rect 265 9 266 17
rect 268 9 269 17
rect 281 9 282 17
rect 284 9 285 17
rect 297 9 298 17
rect 300 9 301 17
rect -10 -44 -9 -36
rect -7 -44 -4 -36
rect 0 -44 3 -36
rect 5 -44 6 -36
rect 18 -44 19 -36
rect 21 -44 22 -36
rect 37 -44 38 -36
rect 40 -44 41 -36
rect 53 -44 54 -36
rect 56 -44 57 -36
rect 69 -44 70 -36
rect 72 -44 73 -36
rect 85 -44 86 -36
rect 88 -44 89 -36
rect 93 -44 94 -36
rect 96 -44 98 -36
rect 102 -44 104 -36
rect 106 -44 107 -36
rect 119 -44 120 -36
rect 122 -44 123 -36
rect 135 -44 136 -36
rect 138 -44 140 -36
rect 144 -44 146 -36
rect 148 -44 149 -36
rect 161 -44 162 -36
rect 164 -44 165 -36
rect 177 -44 178 -36
rect 180 -44 181 -36
rect 185 -44 186 -36
rect 188 -44 189 -36
rect 193 -44 194 -36
rect 196 -44 197 -36
rect 209 -44 210 -36
rect 212 -44 213 -36
rect 225 -44 226 -36
rect 228 -44 234 -36
rect 236 -44 242 -36
rect 244 -44 245 -36
rect 257 -44 258 -36
rect 260 -44 261 -36
rect 273 -44 274 -36
rect 276 -44 277 -36
rect 289 -44 290 -36
rect 292 -44 293 -36
rect 305 -44 306 -36
rect 308 -44 309 -36
rect -10 -97 -9 -89
rect -7 -97 -4 -89
rect 0 -97 3 -89
rect 5 -97 6 -89
rect 18 -97 19 -89
rect 21 -97 22 -89
rect 37 -97 38 -89
rect 40 -97 41 -89
rect 53 -97 54 -89
rect 56 -97 57 -89
rect 69 -97 70 -89
rect 72 -97 73 -89
rect 85 -97 86 -89
rect 88 -97 89 -89
rect 93 -97 94 -89
rect 96 -97 97 -89
rect 101 -97 102 -89
rect 104 -97 106 -89
rect 110 -97 112 -89
rect 114 -97 115 -89
rect 127 -97 128 -89
rect 130 -97 131 -89
rect 143 -97 144 -89
rect 146 -97 147 -89
rect 151 -97 152 -89
rect 154 -97 155 -89
rect 159 -97 160 -89
rect 162 -97 163 -89
rect 167 -97 168 -89
rect 170 -97 171 -89
rect 183 -97 184 -89
rect 186 -97 187 -89
rect 199 -97 200 -89
rect 202 -97 204 -89
rect 208 -97 209 -89
rect 211 -97 212 -89
rect 224 -97 225 -89
rect 227 -97 228 -89
rect 240 -97 241 -89
rect 243 -97 251 -89
rect 253 -97 259 -89
rect 261 -97 267 -89
rect 269 -97 270 -89
rect 282 -97 283 -89
rect 285 -97 286 -89
rect -10 -150 -9 -142
rect -7 -150 -4 -142
rect 0 -150 3 -142
rect 5 -150 6 -142
rect 18 -150 19 -142
rect 21 -150 22 -142
rect 37 -150 38 -142
rect 40 -150 41 -142
rect 53 -150 54 -142
rect 56 -150 57 -142
rect 69 -150 70 -142
rect 72 -150 73 -142
rect 85 -150 86 -142
rect 88 -150 89 -142
rect 93 -150 94 -142
rect 96 -150 97 -142
rect 101 -150 102 -142
rect 104 -150 105 -142
rect 109 -150 110 -142
rect 112 -150 114 -142
rect 118 -150 120 -142
rect 122 -150 123 -142
rect 135 -150 136 -142
rect 138 -150 139 -142
rect 151 -150 152 -142
rect 154 -150 156 -142
rect 160 -150 161 -142
rect 163 -150 164 -142
rect 168 -150 169 -142
rect 171 -150 172 -142
rect 184 -150 185 -142
rect 187 -150 188 -142
rect 200 -150 201 -142
rect 203 -150 205 -142
rect 209 -150 210 -142
rect 212 -150 213 -142
rect 225 -150 226 -142
rect 228 -150 229 -142
rect 241 -150 242 -142
rect 244 -150 250 -142
rect 252 -150 259 -142
rect 261 -150 268 -142
rect 270 -150 277 -142
rect 279 -150 282 -142
rect 294 -150 295 -142
rect 297 -150 298 -142
<< ndcontact >>
rect -14 -15 -10 -11
rect 6 -15 10 -11
rect 14 -15 18 -11
rect 22 -15 26 -11
rect 33 -15 37 -11
rect 41 -15 45 -11
rect 49 -15 53 -11
rect 57 -15 61 -11
rect 65 -15 69 -11
rect 73 -15 77 -11
rect 81 -15 85 -11
rect 89 -15 93 -11
rect 97 -15 101 -11
rect 105 -15 109 -11
rect 113 -15 117 -11
rect 121 -15 125 -11
rect 129 -15 133 -11
rect 147 -15 151 -11
rect 155 -15 159 -11
rect 163 -15 167 -11
rect 171 -15 175 -11
rect 180 -15 184 -11
rect 189 -15 193 -11
rect 197 -15 201 -11
rect 205 -15 209 -11
rect 213 -15 217 -11
rect 221 -15 225 -11
rect 229 -15 233 -11
rect 237 -15 241 -11
rect 245 -15 249 -11
rect 253 -15 257 -11
rect 261 -15 265 -11
rect 269 -15 273 -11
rect 277 -15 281 -11
rect 285 -15 289 -11
rect 293 -15 297 -11
rect 301 -15 305 -11
rect -14 -68 -10 -64
rect 6 -68 10 -64
rect 14 -68 18 -64
rect 22 -68 26 -64
rect 33 -68 37 -64
rect 41 -68 45 -64
rect 49 -68 53 -64
rect 57 -68 61 -64
rect 65 -68 69 -64
rect 73 -68 77 -64
rect 81 -68 85 -64
rect 107 -68 111 -64
rect 115 -68 119 -64
rect 123 -68 127 -64
rect 131 -68 135 -64
rect 149 -68 153 -64
rect 157 -68 161 -64
rect 165 -68 169 -64
rect 173 -68 177 -64
rect 197 -68 201 -64
rect 205 -68 209 -64
rect 213 -68 217 -64
rect 221 -68 225 -64
rect 229 -68 233 -64
rect 237 -68 241 -64
rect 245 -68 249 -64
rect 253 -68 257 -64
rect 261 -68 265 -64
rect 269 -68 273 -64
rect 277 -68 281 -64
rect 285 -68 289 -64
rect 293 -68 297 -64
rect 301 -68 305 -64
rect 309 -68 313 -64
rect -14 -121 -10 -117
rect 6 -121 10 -117
rect 14 -121 18 -117
rect 22 -121 26 -117
rect 33 -121 37 -117
rect 41 -121 45 -117
rect 49 -121 53 -117
rect 57 -121 61 -117
rect 65 -121 69 -117
rect 73 -121 77 -117
rect 81 -121 85 -117
rect 115 -121 119 -117
rect 123 -121 127 -117
rect 131 -121 135 -117
rect 139 -121 143 -117
rect 171 -121 175 -117
rect 179 -121 183 -117
rect 187 -121 191 -117
rect 195 -121 199 -117
rect 212 -121 216 -117
rect 220 -121 224 -117
rect 228 -121 232 -117
rect 236 -121 240 -117
rect 244 -121 248 -117
rect 254 -121 258 -117
rect 262 -121 266 -117
rect 270 -121 274 -117
rect 278 -121 282 -117
rect 286 -121 290 -117
rect -14 -174 -10 -170
rect 6 -174 10 -170
rect 14 -174 18 -170
rect 22 -174 26 -170
rect 33 -174 37 -170
rect 41 -174 45 -170
rect 49 -174 53 -170
rect 57 -174 61 -170
rect 65 -174 69 -170
rect 73 -174 77 -170
rect 81 -174 85 -170
rect 123 -174 127 -170
rect 131 -174 135 -170
rect 139 -174 143 -170
rect 147 -174 151 -170
rect 172 -174 176 -170
rect 180 -174 184 -170
rect 188 -174 192 -170
rect 196 -174 200 -170
rect 213 -174 217 -170
rect 221 -174 225 -170
rect 229 -174 233 -170
rect 237 -174 241 -170
rect 245 -174 249 -170
rect 254 -174 258 -170
rect 263 -174 267 -170
rect 271 -174 275 -170
rect 282 -174 286 -170
rect 290 -174 294 -170
rect 298 -174 302 -170
<< pdcontact >>
rect -14 9 -10 17
rect -4 9 0 17
rect 6 9 10 17
rect 14 9 18 17
rect 22 9 26 17
rect 33 9 37 17
rect 41 9 45 17
rect 49 9 53 17
rect 57 9 61 17
rect 65 9 69 17
rect 73 9 77 17
rect 81 9 85 17
rect 89 9 93 17
rect 97 9 101 17
rect 105 9 109 17
rect 113 9 117 17
rect 121 9 125 17
rect 129 9 133 17
rect 138 9 142 17
rect 147 9 151 17
rect 155 9 159 17
rect 163 9 167 17
rect 171 9 175 17
rect 189 9 193 17
rect 197 9 201 17
rect 205 9 209 17
rect 213 9 217 17
rect 221 9 225 17
rect 229 9 233 17
rect 237 9 241 17
rect 245 9 249 17
rect 253 9 257 17
rect 261 9 265 17
rect 269 9 273 17
rect 277 9 281 17
rect 285 9 289 17
rect 293 9 297 17
rect 301 9 305 17
rect -14 -44 -10 -36
rect -4 -44 0 -36
rect 6 -44 10 -36
rect 14 -44 18 -36
rect 22 -44 26 -36
rect 33 -44 37 -36
rect 41 -44 45 -36
rect 49 -44 53 -36
rect 57 -44 61 -36
rect 65 -44 69 -36
rect 73 -44 77 -36
rect 81 -44 85 -36
rect 89 -44 93 -36
rect 98 -44 102 -36
rect 107 -44 111 -36
rect 115 -44 119 -36
rect 123 -44 127 -36
rect 131 -44 135 -36
rect 140 -44 144 -36
rect 149 -44 153 -36
rect 157 -44 161 -36
rect 165 -44 169 -36
rect 173 -44 177 -36
rect 181 -44 185 -36
rect 189 -44 193 -36
rect 197 -44 201 -36
rect 205 -44 209 -36
rect 213 -44 217 -36
rect 221 -44 225 -36
rect 245 -44 249 -36
rect 253 -44 257 -36
rect 261 -44 265 -36
rect 269 -44 273 -36
rect 277 -44 281 -36
rect 285 -44 289 -36
rect 293 -44 297 -36
rect 301 -44 305 -36
rect 309 -44 313 -36
rect -14 -97 -10 -89
rect -4 -97 0 -89
rect 6 -97 10 -89
rect 14 -97 18 -89
rect 22 -97 26 -89
rect 33 -97 37 -89
rect 41 -97 45 -89
rect 49 -97 53 -89
rect 57 -97 61 -89
rect 65 -97 69 -89
rect 73 -97 77 -89
rect 81 -97 85 -89
rect 89 -97 93 -89
rect 97 -97 101 -89
rect 106 -97 110 -89
rect 115 -97 119 -89
rect 123 -97 127 -89
rect 131 -97 135 -89
rect 139 -97 143 -89
rect 147 -97 151 -89
rect 155 -97 159 -89
rect 163 -97 167 -89
rect 171 -97 175 -89
rect 179 -97 183 -89
rect 187 -97 191 -89
rect 195 -97 199 -89
rect 204 -97 208 -89
rect 212 -97 216 -89
rect 220 -97 224 -89
rect 228 -97 232 -89
rect 236 -97 240 -89
rect 270 -97 274 -89
rect 278 -97 282 -89
rect 286 -97 290 -89
rect -14 -150 -10 -142
rect -4 -150 0 -142
rect 6 -150 10 -142
rect 14 -150 18 -142
rect 22 -150 26 -142
rect 33 -150 37 -142
rect 41 -150 45 -142
rect 49 -150 53 -142
rect 57 -150 61 -142
rect 65 -150 69 -142
rect 73 -150 77 -142
rect 81 -150 85 -142
rect 89 -150 93 -142
rect 97 -150 101 -142
rect 105 -150 109 -142
rect 114 -150 118 -142
rect 123 -150 127 -142
rect 131 -150 135 -142
rect 139 -150 143 -142
rect 147 -150 151 -142
rect 156 -150 160 -142
rect 164 -150 168 -142
rect 172 -150 176 -142
rect 180 -150 184 -142
rect 188 -150 192 -142
rect 196 -150 200 -142
rect 205 -150 209 -142
rect 213 -150 217 -142
rect 221 -150 225 -142
rect 229 -150 233 -142
rect 237 -150 241 -142
rect 282 -150 286 -142
rect 290 -150 294 -142
rect 298 -150 302 -142
<< polysilicon >>
rect -9 17 -7 20
rect 3 17 5 20
rect 19 17 21 20
rect 38 17 40 20
rect 54 17 56 20
rect 70 17 72 27
rect 86 17 88 20
rect 102 17 104 20
rect 118 17 120 27
rect 134 17 136 20
rect 144 17 146 20
rect 160 17 162 20
rect 176 17 178 20
rect 186 17 188 20
rect 202 17 204 20
rect 218 17 220 20
rect 234 17 236 20
rect 250 17 252 23
rect 266 17 268 27
rect 282 17 284 20
rect 298 17 300 27
rect -9 -11 -7 9
rect 3 -11 5 9
rect 19 -11 21 9
rect 38 -11 40 9
rect 54 -11 56 9
rect 70 6 72 9
rect 70 -11 72 -8
rect 86 -11 88 9
rect 102 -11 104 9
rect 118 6 120 9
rect 118 -11 120 -8
rect 134 -11 136 9
rect 144 -11 146 9
rect 160 -11 162 9
rect 176 -11 178 9
rect 186 -11 188 9
rect 202 -11 204 9
rect 218 -11 220 9
rect 234 -11 236 9
rect 250 6 252 9
rect 250 -11 252 -8
rect 266 -11 268 9
rect 282 -11 284 9
rect 298 6 300 9
rect 298 -11 300 -6
rect -9 -18 -7 -15
rect 3 -18 5 -15
rect 19 -18 21 -15
rect 38 -18 40 -15
rect 54 -18 56 -15
rect 70 -22 72 -15
rect -9 -36 -7 -33
rect 3 -36 5 -33
rect 19 -36 21 -33
rect 38 -36 40 -33
rect 54 -36 56 -33
rect 70 -36 72 -26
rect 86 -36 88 -15
rect 102 -27 104 -15
rect 118 -22 120 -15
rect 134 -18 136 -15
rect 144 -18 146 -15
rect 160 -18 162 -15
rect 176 -18 178 -15
rect 94 -29 104 -27
rect 94 -36 96 -29
rect 104 -36 106 -33
rect 120 -36 122 -33
rect 136 -36 138 -33
rect 146 -36 148 -33
rect 162 -36 164 -33
rect 178 -36 180 -33
rect 186 -36 188 -15
rect 202 -18 204 -15
rect 218 -18 220 -15
rect 234 -18 236 -15
rect 250 -22 252 -15
rect 266 -27 268 -15
rect 282 -18 284 -15
rect 298 -22 300 -15
rect 194 -29 268 -27
rect 194 -36 196 -29
rect 210 -36 212 -33
rect 226 -36 228 -33
rect 234 -36 236 -33
rect 242 -36 244 -33
rect 258 -36 260 -33
rect 274 -36 276 -26
rect 290 -36 292 -32
rect 306 -36 308 -26
rect -9 -64 -7 -44
rect 3 -64 5 -44
rect 19 -64 21 -44
rect 38 -64 40 -44
rect 54 -64 56 -44
rect 70 -47 72 -44
rect 70 -64 72 -61
rect 86 -64 88 -44
rect 94 -64 96 -44
rect 104 -64 106 -44
rect 120 -64 122 -44
rect 136 -64 138 -44
rect 146 -64 148 -44
rect 162 -64 164 -44
rect 178 -64 180 -44
rect 186 -64 188 -44
rect 194 -64 196 -44
rect 210 -64 212 -44
rect 226 -64 228 -44
rect 234 -46 236 -44
rect 234 -64 236 -50
rect 242 -64 244 -44
rect 258 -64 260 -44
rect 274 -64 276 -44
rect 290 -64 292 -44
rect 306 -48 308 -44
rect 306 -64 308 -61
rect -9 -71 -7 -68
rect 3 -71 5 -68
rect 19 -71 21 -68
rect 38 -71 40 -68
rect 54 -71 56 -68
rect 70 -75 72 -68
rect -9 -89 -7 -86
rect 3 -89 5 -86
rect 19 -89 21 -86
rect 38 -89 40 -86
rect 54 -89 56 -86
rect 70 -89 72 -79
rect 86 -89 88 -68
rect 94 -89 96 -68
rect 104 -69 106 -68
rect 102 -71 106 -69
rect 120 -71 122 -68
rect 102 -89 104 -71
rect 136 -81 138 -68
rect 146 -76 148 -68
rect 162 -71 164 -68
rect 178 -71 180 -68
rect 186 -71 188 -68
rect 194 -74 196 -68
rect 210 -71 212 -68
rect 226 -71 228 -68
rect 234 -71 236 -68
rect 194 -76 202 -74
rect 242 -76 244 -68
rect 258 -71 260 -68
rect 274 -71 276 -68
rect 290 -73 292 -68
rect 290 -75 294 -73
rect 306 -75 308 -68
rect 146 -78 170 -76
rect 136 -83 162 -81
rect 112 -89 114 -86
rect 128 -89 130 -86
rect 144 -89 146 -86
rect 152 -89 154 -86
rect 160 -89 162 -83
rect 168 -89 170 -78
rect 184 -89 186 -86
rect 200 -89 202 -76
rect 209 -78 244 -76
rect 209 -89 211 -78
rect 225 -89 227 -86
rect 241 -89 243 -86
rect 251 -89 253 -86
rect 259 -89 261 -86
rect 267 -89 269 -86
rect 283 -89 285 -86
rect -9 -117 -7 -97
rect 3 -117 5 -97
rect 19 -117 21 -97
rect 38 -117 40 -97
rect 54 -117 56 -97
rect 70 -100 72 -97
rect 70 -117 72 -114
rect 86 -117 88 -97
rect 94 -117 96 -97
rect 102 -117 104 -97
rect 112 -117 114 -97
rect 128 -117 130 -97
rect 144 -117 146 -97
rect 152 -106 154 -97
rect 152 -117 154 -110
rect 160 -117 162 -97
rect 168 -117 170 -97
rect 184 -117 186 -97
rect 200 -117 202 -97
rect 209 -106 211 -97
rect 210 -110 211 -106
rect 209 -117 211 -110
rect 225 -117 227 -97
rect 241 -117 243 -97
rect 251 -104 253 -97
rect 259 -104 261 -97
rect 252 -108 253 -104
rect 251 -117 253 -108
rect 259 -117 261 -108
rect 267 -117 269 -97
rect 283 -117 285 -97
rect -9 -124 -7 -121
rect 3 -124 5 -121
rect 19 -124 21 -121
rect 38 -124 40 -121
rect 54 -124 56 -121
rect 70 -128 72 -121
rect -9 -142 -7 -139
rect 3 -142 5 -139
rect 19 -142 21 -139
rect 38 -142 40 -139
rect 54 -142 56 -139
rect 70 -142 72 -132
rect 86 -142 88 -121
rect 94 -142 96 -121
rect 102 -142 104 -121
rect 112 -122 114 -121
rect 110 -124 114 -122
rect 128 -124 130 -121
rect 110 -142 112 -124
rect 144 -130 146 -121
rect 120 -132 146 -130
rect 152 -130 154 -121
rect 160 -124 162 -121
rect 168 -124 170 -121
rect 184 -124 186 -121
rect 200 -124 202 -121
rect 209 -124 211 -121
rect 225 -124 227 -121
rect 241 -124 243 -121
rect 251 -124 253 -121
rect 259 -124 261 -121
rect 267 -129 269 -121
rect 283 -124 285 -121
rect 292 -129 294 -75
rect 152 -132 171 -130
rect 120 -142 122 -132
rect 136 -142 138 -139
rect 152 -142 154 -139
rect 161 -142 163 -139
rect 169 -142 171 -132
rect 201 -131 269 -129
rect 284 -131 294 -129
rect 185 -142 187 -139
rect 201 -142 203 -131
rect 284 -134 286 -131
rect 210 -136 286 -134
rect 210 -142 212 -136
rect 226 -142 228 -139
rect 242 -142 244 -139
rect 250 -142 252 -139
rect 259 -142 261 -139
rect 268 -142 270 -139
rect 277 -142 279 -139
rect 295 -142 297 -139
rect -9 -170 -7 -150
rect 3 -170 5 -150
rect 19 -170 21 -150
rect 38 -170 40 -150
rect 54 -170 56 -150
rect 70 -153 72 -150
rect 70 -170 72 -167
rect 86 -170 88 -150
rect 94 -170 96 -150
rect 102 -170 104 -150
rect 110 -170 112 -150
rect 120 -170 122 -150
rect 136 -170 138 -150
rect 152 -170 154 -150
rect 161 -165 163 -150
rect 162 -169 163 -165
rect 161 -170 163 -169
rect 169 -170 171 -150
rect 185 -170 187 -150
rect 201 -157 203 -150
rect 202 -161 203 -157
rect 210 -159 212 -150
rect 201 -170 203 -161
rect 211 -163 212 -159
rect 210 -170 212 -163
rect 226 -170 228 -150
rect 242 -170 244 -150
rect 250 -157 252 -150
rect 259 -157 261 -150
rect 268 -157 270 -150
rect 277 -157 279 -150
rect 250 -170 252 -161
rect 259 -170 261 -161
rect 268 -170 270 -161
rect 277 -170 279 -161
rect 295 -170 297 -150
rect -9 -177 -7 -174
rect 3 -177 5 -174
rect 19 -177 21 -174
rect 38 -177 40 -174
rect 54 -177 56 -174
rect 70 -181 72 -174
rect 86 -177 88 -174
rect 94 -177 96 -174
rect 102 -177 104 -174
rect 110 -177 112 -174
rect 120 -177 122 -174
rect 136 -177 138 -174
rect 152 -177 154 -174
rect 161 -177 163 -174
rect 169 -177 171 -174
rect 185 -177 187 -174
rect 201 -177 203 -174
rect 210 -177 212 -174
rect 226 -177 228 -174
rect 242 -177 244 -174
rect 250 -177 252 -174
rect 259 -177 261 -174
rect 268 -177 270 -174
rect 277 -177 279 -174
rect 295 -177 297 -174
<< polycontact >>
rect 66 23 70 27
rect 114 23 118 27
rect 248 23 252 27
rect 268 23 272 27
rect 294 23 298 27
rect -13 -1 -9 3
rect -1 -10 3 -6
rect 15 -2 19 2
rect 34 -1 38 3
rect 50 -1 54 3
rect 82 -8 86 -4
rect 98 -2 102 2
rect 130 -3 134 1
rect 140 -4 144 0
rect 156 -2 160 2
rect 172 -1 176 3
rect 182 -2 186 2
rect 198 -2 202 2
rect 214 -2 218 2
rect 230 -1 234 3
rect 278 -1 282 3
rect 66 -22 70 -18
rect 66 -30 70 -26
rect 114 -22 118 -18
rect 246 -22 250 -18
rect 294 -22 298 -18
rect 276 -30 280 -26
rect 302 -30 306 -26
rect -13 -54 -9 -50
rect -1 -63 3 -59
rect 15 -55 19 -51
rect 34 -54 38 -50
rect 50 -54 54 -50
rect 100 -57 104 -53
rect 116 -55 120 -51
rect 132 -55 136 -51
rect 142 -63 146 -59
rect 158 -55 162 -51
rect 174 -55 178 -51
rect 206 -55 210 -51
rect 222 -57 226 -53
rect 232 -50 236 -46
rect 254 -56 258 -52
rect 270 -55 274 -51
rect 286 -55 290 -51
rect 66 -75 70 -71
rect 66 -83 70 -79
rect 302 -75 306 -71
rect -13 -107 -9 -103
rect -1 -116 3 -112
rect 15 -108 19 -104
rect 34 -107 38 -103
rect 50 -107 54 -103
rect 108 -110 112 -106
rect 124 -108 128 -104
rect 150 -110 154 -106
rect 180 -108 184 -104
rect 196 -108 200 -104
rect 206 -110 210 -106
rect 221 -108 225 -104
rect 237 -108 241 -104
rect 248 -108 252 -104
rect 257 -108 261 -104
rect 279 -108 283 -104
rect 66 -128 70 -124
rect 66 -136 70 -132
rect -13 -160 -9 -156
rect -1 -169 3 -165
rect 15 -161 19 -157
rect 34 -160 38 -156
rect 50 -160 54 -156
rect 116 -163 120 -159
rect 132 -161 136 -157
rect 148 -161 152 -157
rect 158 -169 162 -165
rect 181 -161 185 -157
rect 198 -161 202 -157
rect 207 -163 211 -159
rect 222 -161 226 -157
rect 238 -161 242 -157
rect 248 -161 252 -157
rect 257 -161 261 -157
rect 266 -161 270 -157
rect 275 -161 279 -157
rect 291 -161 295 -157
rect 66 -181 70 -177
<< metal1 >>
rect -20 23 -2 26
rect -14 17 -10 23
rect 3 23 20 26
rect 25 23 37 26
rect 6 17 10 23
rect 14 17 18 23
rect 33 17 37 23
rect 134 23 204 27
rect 49 17 53 22
rect 81 17 85 22
rect 97 17 101 22
rect 129 17 133 23
rect 147 17 151 23
rect -4 6 0 9
rect -4 3 10 6
rect 6 2 10 3
rect 6 -2 15 2
rect 6 -11 10 -2
rect 22 -11 26 9
rect 41 -11 45 9
rect 57 -11 61 9
rect 65 3 69 9
rect 66 -2 69 3
rect -14 -19 -10 -15
rect 14 -18 18 -15
rect -20 -22 10 -19
rect 15 -22 18 -18
rect 65 -11 69 -2
rect 73 -5 77 9
rect 82 -4 86 -1
rect 73 -11 77 -10
rect 89 -11 93 9
rect 105 2 109 9
rect 113 2 117 9
rect 98 -3 102 -2
rect 105 -2 117 2
rect 105 -11 109 -2
rect 113 -11 117 -2
rect 155 17 159 23
rect 171 17 175 23
rect 197 17 201 23
rect 209 23 217 27
rect 213 17 217 23
rect 272 23 294 27
rect 229 17 233 22
rect 261 17 265 22
rect 277 17 281 23
rect 121 -3 125 9
rect 138 6 142 9
rect 138 3 151 6
rect 147 2 151 3
rect 163 3 167 9
rect 121 -11 125 -8
rect 147 -2 156 2
rect 163 -1 172 3
rect 147 -11 151 -2
rect 163 -11 167 -1
rect 189 2 193 9
rect 205 2 209 9
rect 189 -2 198 2
rect 205 -2 214 2
rect 189 -5 193 -2
rect 180 -8 193 -5
rect 180 -11 184 -8
rect 205 -11 209 -2
rect 221 -11 225 9
rect 237 3 241 9
rect 245 3 249 9
rect 237 -2 249 3
rect 237 -11 241 -2
rect 33 -19 37 -15
rect 49 -19 53 -15
rect 81 -18 85 -15
rect 33 -22 45 -19
rect 49 -22 66 -19
rect 73 -22 85 -18
rect 97 -19 101 -15
rect 97 -22 114 -19
rect 129 -19 133 -15
rect 155 -19 159 -15
rect 171 -19 175 -15
rect 189 -18 193 -15
rect 245 -11 249 -2
rect 253 -1 257 9
rect 253 -11 257 -6
rect 269 -11 273 9
rect 285 3 289 9
rect 293 3 297 9
rect 285 -2 297 3
rect 285 -11 289 -2
rect 293 -11 297 -2
rect 301 -5 305 9
rect 301 -11 305 -10
rect 197 -18 201 -15
rect 213 -18 217 -15
rect 189 -19 201 -18
rect 212 -19 217 -18
rect 229 -19 233 -15
rect 261 -18 265 -15
rect 127 -22 225 -19
rect 229 -22 246 -19
rect 260 -22 265 -18
rect 277 -19 281 -15
rect 277 -22 294 -19
rect -20 -30 -2 -27
rect -14 -36 -10 -30
rect 3 -30 37 -27
rect 6 -36 10 -30
rect 14 -36 18 -30
rect 33 -36 37 -30
rect 158 -28 176 -25
rect 81 -31 128 -28
rect 49 -36 53 -31
rect 81 -36 85 -31
rect 98 -32 128 -31
rect 98 -36 102 -32
rect 115 -36 119 -32
rect 133 -32 161 -28
rect 173 -31 273 -28
rect 280 -30 302 -26
rect 133 -33 135 -32
rect 131 -36 135 -33
rect 149 -36 153 -32
rect -4 -47 0 -44
rect -4 -50 10 -47
rect 6 -51 10 -50
rect 6 -55 15 -51
rect 6 -64 10 -55
rect 22 -64 26 -44
rect 41 -64 45 -44
rect 57 -64 61 -44
rect 65 -50 69 -44
rect 66 -55 69 -50
rect -14 -72 -10 -68
rect 14 -71 18 -68
rect -20 -75 10 -72
rect 15 -75 18 -71
rect 65 -64 69 -55
rect 157 -36 161 -32
rect 173 -36 177 -31
rect 189 -36 193 -31
rect 205 -36 209 -31
rect 221 -36 225 -31
rect 253 -36 257 -31
rect 269 -36 273 -31
rect 285 -36 289 -30
rect 73 -58 77 -44
rect 89 -47 93 -44
rect 107 -47 111 -44
rect 89 -50 111 -47
rect 107 -51 111 -50
rect 123 -46 127 -44
rect 140 -47 144 -44
rect 140 -50 153 -47
rect 149 -51 153 -50
rect 100 -58 104 -57
rect 107 -55 116 -51
rect 73 -64 77 -63
rect 107 -64 111 -55
rect 123 -64 127 -51
rect 149 -55 158 -51
rect 149 -64 153 -55
rect 165 -64 169 -44
rect 181 -47 185 -44
rect 197 -47 201 -44
rect 181 -50 201 -47
rect 197 -51 201 -50
rect 197 -55 206 -51
rect 197 -64 201 -55
rect 213 -58 217 -44
rect 245 -52 249 -44
rect 261 -46 265 -44
rect 245 -56 254 -52
rect 245 -58 249 -56
rect 229 -61 249 -58
rect 213 -64 217 -63
rect 229 -64 233 -61
rect 245 -64 249 -61
rect 261 -64 265 -51
rect 277 -64 281 -44
rect 293 -51 297 -44
rect 301 -51 305 -44
rect 293 -55 305 -51
rect 293 -64 297 -55
rect 301 -64 305 -55
rect 309 -55 313 -44
rect 309 -64 313 -60
rect 33 -72 37 -68
rect 49 -72 53 -68
rect 33 -75 45 -72
rect 49 -75 66 -72
rect 81 -72 85 -68
rect 115 -72 119 -68
rect 131 -72 135 -68
rect 157 -72 161 -68
rect 173 -72 177 -68
rect 205 -72 209 -68
rect 221 -72 225 -68
rect 237 -72 241 -68
rect 253 -72 257 -68
rect 269 -72 273 -68
rect 80 -75 273 -72
rect 285 -72 289 -68
rect 285 -75 302 -72
rect -20 -83 -2 -80
rect -14 -89 -10 -83
rect 3 -83 37 -80
rect 6 -89 10 -83
rect 14 -89 18 -83
rect 33 -89 37 -83
rect 181 -80 198 -78
rect 81 -81 300 -80
rect 81 -83 184 -81
rect 195 -83 300 -81
rect 49 -89 53 -84
rect 81 -89 85 -83
rect 97 -89 101 -83
rect 115 -89 119 -83
rect -4 -100 0 -97
rect -4 -103 10 -100
rect 6 -104 10 -103
rect 6 -108 15 -104
rect 6 -117 10 -108
rect 22 -117 26 -97
rect 41 -117 45 -97
rect 57 -117 61 -97
rect 65 -103 69 -97
rect 66 -108 69 -103
rect -14 -125 -10 -121
rect 14 -124 18 -121
rect -20 -128 10 -125
rect 15 -128 18 -124
rect 65 -117 69 -108
rect 123 -89 127 -83
rect 139 -89 143 -83
rect 163 -89 167 -83
rect 179 -89 183 -83
rect 195 -89 199 -83
rect 212 -89 216 -83
rect 220 -89 224 -83
rect 236 -89 240 -83
rect 278 -89 282 -83
rect 73 -111 77 -97
rect 89 -100 93 -97
rect 106 -100 110 -97
rect 131 -99 135 -97
rect 89 -103 119 -100
rect 115 -104 119 -103
rect 155 -100 159 -97
rect 171 -100 175 -97
rect 155 -103 175 -100
rect 171 -104 175 -103
rect 115 -108 124 -104
rect 73 -117 77 -116
rect 115 -117 119 -108
rect 131 -117 135 -104
rect 171 -108 180 -104
rect 171 -117 175 -108
rect 187 -117 191 -97
rect 204 -100 208 -97
rect 204 -103 216 -100
rect 213 -104 216 -103
rect 228 -104 232 -97
rect 213 -108 221 -104
rect 228 -108 237 -104
rect 245 -108 248 -101
rect 270 -104 274 -97
rect 270 -108 279 -104
rect 213 -117 216 -108
rect 228 -117 232 -108
rect 270 -111 274 -108
rect 244 -114 274 -111
rect 244 -117 248 -114
rect 262 -117 266 -114
rect 286 -117 290 -102
rect 33 -125 37 -121
rect 49 -125 53 -121
rect 33 -128 45 -125
rect 49 -128 66 -125
rect 81 -125 85 -121
rect 123 -125 127 -121
rect 139 -125 143 -121
rect 179 -125 183 -121
rect 195 -125 199 -121
rect 220 -125 224 -121
rect 236 -125 240 -121
rect 254 -125 258 -121
rect 270 -125 274 -121
rect 278 -125 282 -121
rect 81 -128 287 -125
rect -20 -136 -2 -133
rect -14 -142 -10 -136
rect 3 -136 37 -133
rect 6 -142 10 -136
rect 14 -142 18 -136
rect 33 -142 37 -136
rect 297 -133 300 -83
rect 81 -136 300 -133
rect 49 -142 53 -137
rect 81 -142 85 -136
rect 97 -142 101 -136
rect 114 -142 118 -136
rect 131 -142 135 -136
rect 147 -142 151 -136
rect 164 -142 168 -136
rect 180 -142 184 -136
rect 196 -142 200 -136
rect 213 -142 217 -136
rect -4 -153 0 -150
rect -4 -156 10 -153
rect 6 -157 10 -156
rect 6 -161 15 -157
rect 6 -170 10 -161
rect 22 -170 26 -150
rect 41 -170 45 -150
rect 57 -170 61 -150
rect 65 -156 69 -150
rect 66 -161 69 -156
rect -14 -178 -10 -174
rect 14 -178 18 -174
rect -20 -182 10 -178
rect 15 -183 18 -178
rect 65 -170 69 -161
rect 221 -142 225 -136
rect 237 -142 241 -136
rect 290 -142 294 -136
rect 73 -164 77 -150
rect 89 -153 93 -150
rect 105 -153 109 -150
rect 123 -153 127 -150
rect 89 -156 127 -153
rect 123 -157 127 -156
rect 139 -152 143 -150
rect 156 -153 160 -150
rect 172 -153 176 -150
rect 156 -156 176 -153
rect 172 -157 176 -156
rect 188 -152 192 -150
rect 205 -153 209 -150
rect 205 -156 217 -153
rect 214 -157 217 -156
rect 229 -157 233 -150
rect 123 -161 132 -157
rect 73 -170 77 -169
rect 123 -170 127 -161
rect 139 -170 143 -157
rect 172 -161 181 -157
rect 172 -170 176 -161
rect 188 -170 192 -157
rect 214 -161 222 -157
rect 229 -161 238 -157
rect 282 -157 286 -150
rect 282 -161 291 -157
rect 214 -170 217 -161
rect 229 -170 233 -161
rect 282 -164 286 -161
rect 245 -167 286 -164
rect 245 -170 249 -167
rect 263 -170 267 -167
rect 282 -170 286 -167
rect 298 -170 302 -150
rect 33 -178 37 -174
rect 49 -178 53 -174
rect 33 -181 45 -178
rect 49 -181 66 -178
rect 81 -178 85 -174
rect 131 -178 135 -174
rect 147 -178 151 -174
rect 180 -178 184 -174
rect 196 -178 200 -174
rect 221 -178 225 -174
rect 237 -178 241 -174
rect 254 -178 258 -174
rect 271 -178 275 -174
rect 290 -178 294 -174
rect 81 -181 302 -178
rect 37 -182 45 -181
<< m2contact >>
rect 49 22 54 27
rect 61 22 66 27
rect 96 22 101 27
rect 109 22 114 27
rect -18 -2 -13 3
rect -6 -10 -1 -5
rect 29 -2 34 3
rect 49 -6 54 -1
rect 61 -2 66 3
rect 81 -1 86 4
rect 72 -10 77 -5
rect 97 -8 102 -3
rect 228 22 233 27
rect 243 22 248 27
rect 129 1 134 6
rect 120 -8 125 -3
rect 139 -9 144 -4
rect 181 2 186 7
rect 213 -7 218 -2
rect 22 -20 27 -15
rect 277 -6 282 -1
rect 301 -10 306 -5
rect 49 -31 54 -26
rect 61 -31 66 -26
rect -18 -55 -13 -50
rect -6 -63 -1 -58
rect 29 -55 34 -50
rect 49 -59 54 -54
rect 165 -36 170 -31
rect 72 -63 77 -58
rect 141 -59 146 -54
rect 230 -55 235 -50
rect 261 -51 266 -46
rect 213 -63 218 -58
rect 269 -60 274 -55
rect 285 -60 290 -55
rect 309 -60 314 -55
rect 22 -73 27 -68
rect 49 -84 54 -79
rect 61 -84 66 -79
rect -18 -108 -13 -103
rect -6 -116 -1 -111
rect 29 -108 34 -103
rect 49 -112 54 -107
rect 131 -104 136 -99
rect 72 -116 77 -111
rect 244 -101 249 -96
rect 255 -104 260 -99
rect 286 -102 291 -97
rect 204 -115 209 -110
rect 22 -126 27 -121
rect 49 -137 54 -132
rect 61 -137 66 -132
rect -18 -161 -13 -156
rect -6 -169 -1 -164
rect 29 -161 34 -156
rect 49 -165 54 -160
rect 188 -157 193 -152
rect 246 -157 252 -151
rect 72 -169 77 -164
rect 156 -165 161 -160
rect 196 -166 201 -161
rect 32 -186 37 -181
<< metal2 >>
rect 29 23 49 26
rect 29 3 32 23
rect 54 23 61 27
rect 89 23 96 27
rect 89 4 92 23
rect 101 23 109 27
rect -13 -1 29 3
rect 66 -1 81 3
rect 86 -1 92 4
rect 105 6 109 23
rect 213 23 228 27
rect 105 3 129 6
rect 168 3 181 7
rect -1 -10 72 -6
rect 102 -8 120 -4
rect 125 -9 139 -5
rect 168 -15 171 3
rect 213 -2 216 23
rect 233 23 243 27
rect 27 -18 171 -15
rect 277 -10 301 -6
rect 54 -30 61 -26
rect 29 -34 54 -31
rect 29 -50 32 -34
rect -13 -54 29 -50
rect 142 -54 146 -18
rect 277 -27 282 -10
rect 261 -30 282 -27
rect 170 -36 235 -33
rect 231 -50 235 -36
rect -1 -63 72 -59
rect 261 -46 265 -30
rect 290 -60 309 -57
rect 27 -71 91 -68
rect 54 -83 61 -79
rect 29 -87 54 -84
rect 29 -103 32 -87
rect -13 -107 29 -103
rect -1 -116 72 -112
rect 27 -124 84 -121
rect 54 -136 61 -132
rect 29 -140 54 -137
rect 29 -156 32 -140
rect -13 -160 29 -156
rect -1 -169 72 -165
rect 81 -175 84 -124
rect 88 -122 91 -71
rect 213 -80 216 -63
rect 270 -76 274 -60
rect 270 -79 289 -76
rect 213 -83 249 -80
rect 245 -96 249 -83
rect 136 -103 220 -100
rect 286 -97 289 -79
rect 204 -122 209 -115
rect 88 -125 209 -122
rect 217 -122 220 -103
rect 255 -122 258 -104
rect 217 -125 258 -122
rect 164 -129 168 -125
rect 156 -132 168 -129
rect 156 -160 160 -132
rect 193 -157 246 -154
rect 196 -175 200 -166
rect 81 -178 200 -175
rect 10 -186 32 -183
<< m123contact >>
rect -2 22 3 27
rect 20 23 25 28
rect 80 22 85 27
rect 129 23 134 28
rect 204 22 209 27
rect 260 22 265 27
rect 229 -6 234 -1
rect 253 -6 258 -1
rect 10 -23 15 -18
rect -2 -31 3 -26
rect 40 -27 45 -22
rect 73 -27 78 -22
rect 128 -33 133 -28
rect 61 -55 66 -50
rect 123 -51 128 -46
rect 221 -53 226 -48
rect 99 -63 104 -58
rect 131 -60 136 -55
rect 173 -60 178 -55
rect 10 -76 15 -71
rect -2 -84 3 -79
rect 40 -80 45 -75
rect 61 -108 66 -103
rect 10 -129 15 -124
rect -2 -137 3 -132
rect 40 -133 45 -128
rect 61 -161 66 -156
rect 10 -183 15 -178
rect 22 -179 27 -174
rect 187 -89 192 -84
rect 107 -115 112 -110
rect 149 -115 154 -110
rect 195 -113 200 -108
rect 139 -157 144 -152
rect 256 -157 261 -152
rect 265 -157 270 -152
rect 274 -157 279 -152
rect 115 -168 120 -163
rect 147 -166 152 -161
rect 205 -168 210 -163
<< metal3 >>
rect 25 23 80 26
rect 0 -26 3 22
rect 41 -22 76 -19
rect 0 -79 3 -31
rect 11 -71 14 -23
rect 41 -75 45 -27
rect 129 -28 133 23
rect 209 23 260 27
rect 234 -6 253 -3
rect 229 -24 234 -6
rect 229 -27 242 -24
rect 128 -48 226 -46
rect 128 -50 221 -48
rect 66 -55 93 -52
rect 90 -59 93 -55
rect 90 -63 99 -59
rect 104 -60 131 -59
rect 136 -60 173 -56
rect 238 -58 242 -27
rect 178 -60 242 -58
rect 104 -63 136 -60
rect 173 -62 242 -60
rect 0 -132 3 -84
rect 11 -124 14 -76
rect 41 -128 45 -80
rect 192 -89 285 -85
rect 66 -108 92 -104
rect 89 -112 92 -108
rect 89 -115 107 -112
rect 112 -113 149 -110
rect 154 -113 195 -110
rect 282 -125 285 -89
rect 11 -132 40 -129
rect 11 -178 14 -132
rect 274 -128 285 -125
rect 234 -136 268 -133
rect 234 -153 237 -136
rect 265 -152 268 -136
rect 274 -152 277 -128
rect 144 -156 237 -153
rect 66 -161 100 -158
rect 97 -164 100 -161
rect 97 -167 115 -164
rect 120 -166 147 -163
rect 152 -166 205 -163
rect 256 -176 259 -157
rect 27 -179 259 -176
<< labels >>
rlabel m2contact -16 0 -16 0 3 A0
rlabel m2contact -4 -8 -4 -8 1 B0
rlabel metal1 8 -4 8 -4 1 D0
rlabel metal1 24 -3 24 -3 1 G0
rlabel m2contact 63 0 63 0 1 P0
rlabel m2contact -16 -53 -16 -53 3 A1
rlabel m2contact -4 -61 -4 -61 1 B1
rlabel metal1 8 -57 8 -57 1 D1
rlabel metal1 24 -56 24 -56 1 G1
rlabel metal1 -13 25 -13 25 5 vdd
rlabel metal1 -13 -21 -13 -21 1 gnd
rlabel m123contact 63 -160 63 -160 1 P3
rlabel metal1 24 -110 24 -110 1 G2
rlabel metal1 24 -163 24 -163 1 G3
rlabel metal1 8 -110 8 -110 1 D2
rlabel metal1 7 -163 7 -163 1 D3
rlabel m2contact -3 -167 -3 -167 1 B3
rlabel m2contact -16 -160 -16 -160 3 A3
rlabel m2contact -4 -114 -4 -114 1 B2
rlabel m2contact -16 -107 -16 -107 3 A2
rlabel m2contact 99 -5 99 -5 1 C0
rlabel metal1 111 0 111 0 1 S0
rlabel metal1 207 -1 207 -1 1 C1
rlabel metal1 164 0 164 0 1 E1
rlabel m123contact 63 -52 63 -52 1 P1
rlabel metal1 125 -58 125 -58 1 E3
rlabel metal1 167 -55 167 -55 1 E2
rlabel metal1 133 -107 133 -107 1 E6
rlabel metal1 63 -106 63 -105 1 P2
rlabel metal1 141 -161 141 -161 1 E10
rlabel metal1 190 -159 190 -159 1 E8
rlabel metal1 231 -161 231 -161 1 E7
rlabel metal1 215 -53 215 -53 1 E5
rlabel metal1 291 0 291 0 1 S2
rlabel metal1 299 -53 299 -53 1 S3
rlabel metal1 300 -161 300 -161 1 C4
rlabel metal1 243 0 243 0 1 S1
rlabel metal1 262 -56 262 -56 1 C2
rlabel metal1 142 26 142 26 5 vdd
rlabel metal1 139 -21 139 -21 1 gnd
rlabel metal1 113 -30 113 -30 1 vdd
rlabel metal1 262 -20 262 -20 1 gnd
rlabel metal1 263 -74 263 -74 1 gnd
rlabel metal1 277 -179 277 -179 1 gnd
rlabel metal1 111 -81 111 -81 1 vdd
rlabel metal1 189 -108 189 -108 1 E9
rlabel metal1 230 -106 230 -106 1 E4
rlabel metal1 288 -108 288 -108 1 C3
rlabel metal1 271 -127 271 -127 1 gnd
<< end >>
